`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/26/2018 11:21:36 AM
// Design Name: 
// Module Name: block_classify
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module block_classify(
    input [127:0] input_block,
    input [127:0] bg_block,
    output [127:0] bin_block
    );
endmodule
